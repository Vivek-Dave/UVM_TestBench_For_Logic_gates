
interface intf(input bit clk);
    // ------------------- port declaration-------------------------------------
    logic a;
    logic b;
    
    logic andd;
    logic orr;
    logic nott_a;
    logic nott_b;
    logic xorr;
    logic xnorr;
    logic buff_a;
    logic buff_b;
    logic nandd;
    logic norr;
  	logic temp;
    //--------------------------------------------------------------------------
    //--------------------------------------------------------------------------
        
endinterface

